library ieee;
use ieee.std_logic_1164.all;

----------------------------------------------------------------------
entity adder16 is
	port (
		a		: in  std_logic_vector(15 downto 0);
		b		: in  std_logic_vector(15 downto 0);
		c_in		: in  std_logic;
		sum		: out std_logic_vector(15 downto 0)
	);
end adder16;
----------------------------------------------------------------------

----------------------------------------------------------------------
architecture struct of adder16 is
	signal p, g		: std_logic_vector(15 downto 0);
	signal carry		: std_logic_vector(15 downto 0);
	signal p2, g2		: std_logic_vector(2 downto 0);
	signal carry2		: std_logic_vector(3 downto 0);
	signal net_0		: std_logic;
	signal net_1		: std_logic;
	signal net_2		: std_logic;
	signal net_3		: std_logic;
	signal net_4		: std_logic;
	signal net_5		: std_logic;
	signal net_6		: std_logic;
	signal net_7		: std_logic;
	signal net_8		: std_logic;
	signal net_9		: std_logic;
	signal net_10		: std_logic;
	signal net_11		: std_logic;
	signal net_12		: std_logic;
	signal net_13		: std_logic;
	signal net_14		: std_logic;
	signal net_15		: std_logic;
	signal net_16		: std_logic;
	signal net_17		: std_logic;
	signal net_18		: std_logic;
	signal net_19		: std_logic;
	signal net_20		: std_logic;
	signal net_21		: std_logic;
	signal net_22		: std_logic;
	signal net_23		: std_logic;
	signal net_24		: std_logic;
	signal net_25		: std_logic;
	signal net_26		: std_logic;
	signal net_27		: std_logic;
	signal net_28		: std_logic;
	signal net_29		: std_logic;
	signal net_30		: std_logic;
	signal net_31		: std_logic;
	signal net_32		: std_logic;
	signal net_33		: std_logic;
	signal net_34		: std_logic;
	signal net_35		: std_logic;
	signal net_36		: std_logic;
	signal net_37		: std_logic;
	signal net_38		: std_logic;
begin
	carry(0) <= c_in;
	U1 : XOR2 port map (A1 => a(0), A2 => b(0), Z => p(0));
	U2 : AND2 port map (A1 => a(0), A2 => b(0), Z => g(0));
	U3 : XOR2 port map (A1 => a(1), A2 => b(1), Z => p(1));
	U4 : AND2 port map (A1 => a(1), A2 => b(1), Z => g(1));
	U5 : XOR2 port map (A1 => a(2), A2 => b(2), Z => p(2));
	U6 : AND2 port map (A1 => a(2), A2 => b(2), Z => g(2));
	U7 : XOR2 port map (A1 => a(3), A2 => b(3), Z => p(3));
	U8 : AND2 port map (A1 => a(3), A2 => b(3), Z => g(3));
	U9 : XOR2 port map (A1 => a(4), A2 => b(4), Z => p(4));
	U10 : AND2 port map (A1 => a(4), A2 => b(4), Z => g(4));
	U11 : XOR2 port map (A1 => a(5), A2 => b(5), Z => p(5));
	U12 : AND2 port map (A1 => a(5), A2 => b(5), Z => g(5));
	U13 : XOR2 port map (A1 => a(6), A2 => b(6), Z => p(6));
	U14 : AND2 port map (A1 => a(6), A2 => b(6), Z => g(6));
	U15 : XOR2 port map (A1 => a(7), A2 => b(7), Z => p(7));
	U16 : AND2 port map (A1 => a(7), A2 => b(7), Z => g(7));
	U17 : XOR2 port map (A1 => a(8), A2 => b(8), Z => p(8));
	U18 : AND2 port map (A1 => a(8), A2 => b(8), Z => g(8));
	U19 : XOR2 port map (A1 => a(9), A2 => b(9), Z => p(9));
	U20 : AND2 port map (A1 => a(9), A2 => b(9), Z => g(9));
	U21 : XOR2 port map (A1 => a(10), A2 => b(10), Z => p(10));
	U22 : AND2 port map (A1 => a(10), A2 => b(10), Z => g(10));
	U23 : XOR2 port map (A1 => a(11), A2 => b(11), Z => p(11));
	U24 : AND2 port map (A1 => a(11), A2 => b(11), Z => g(11));
	U25 : XOR2 port map (A1 => a(12), A2 => b(12), Z => p(12));
	U26 : AND2 port map (A1 => a(12), A2 => b(12), Z => g(12));
	U27 : XOR2 port map (A1 => a(13), A2 => b(13), Z => p(13));
	U28 : AND2 port map (A1 => a(13), A2 => b(13), Z => g(13));
	U29 : XOR2 port map (A1 => a(14), A2 => b(14), Z => p(14));
	U30 : AND2 port map (A1 => a(14), A2 => b(14), Z => g(14));
	U31 : XOR2 port map (A1 => a(15), A2 => b(15), Z => p(15));
	U32 : AND2 port map (A1 => a(15), A2 => b(15), Z => g(15));
	U33 : AND4 port map (A1 => p(0), A2 => p(1), A3 => p(2), A4 => p(3), Z => p2(0));
	U34 : AND4 port map (A1 => p(4), A2 => p(5), A3 => p(6), A4 => p(7), Z => p2(1));
	U35 : AND4 port map (A1 => p(8), A2 => p(9), A3 => p(10), A4 => p(11), Z => p2(2));
	U36 : AND4 port map (A1 => g(0), A2 => p(1), A3 => p(2), A4 => p(3), Z => net_0);
	U37 : AND3 port map (A1 => g(1), A2 => p(2), A3 => p(3), Z => net_1);
	U38 : AND2 port map (A1 => g(2), A2 => p(3), Z => net_2);
	U39 : OR4 port map (A1 => net_0, A2 => net_1, A3 => net_2, A4 => g(3), Z => g2(0));
	U40 : AND4 port map (A1 => g(4), A2 => p(5), A3 => p(6), A4 => p(7), Z => net_3);
	U41 : AND3 port map (A1 => g(5), A2 => p(6), A3 => p(7), Z => net_4);
	U42 : AND2 port map (A1 => g(6), A2 => p(7), Z => net_5);
	U43 : OR4 port map (A1 => net_3, A2 => net_4, A3 => net_5, A4 => g(7), Z => g2(1));
	U44 : AND4 port map (A1 => g(8), A2 => p(9), A3 => p(10), A4 => p(11), Z => net_6);
	U45 : AND3 port map (A1 => g(9), A2 => p(10), A3 => p(11), Z => net_7);
	U46 : AND2 port map (A1 => g(10), A2 => p(11), Z => net_8);
	U47 : OR4 port map (A1 => net_6, A2 => net_7, A3 => net_8, A4 => g(11), Z => g2(2));
	carry2(0) <= carry(0);
	U48 : AND4 port map (A1 => carry2(0), A2 => p2(0), A3 => p2(1), A4 => p2(2), Z => net_9);
	U49 : AND3 port map (A1 => g2(0), A2 => p2(1), A3 => p2(2), Z => net_10);
	U50 : AND2 port map (A1 => g2(1), A2 => p2(2), Z => net_11);
	U51 : OR4 port map (A1 => net_9, A2 => net_10, A3 => net_11, A4 => g2(2), Z => carry2(3));
	U52 : AND3 port map (A1 => carry2(0), A2 => p2(0), A3 => p2(1), Z => net_12);
	U53 : AND2 port map (A1 => g2(0), A2 => p2(1), Z => net_13);
	U54 : OR3 port map (A1 => net_12, A2 => net_13, A3 => g2(1), Z => carry2(2));
	U55 : AND2 port map (A1 => carry2(0), A2 => p2(0), Z => net_14);
	U56 : OR2 port map (A1 => net_14, A2 => g2(0), Z => carry2(1));
	U57 : AND4 port map (A1 => carry(0), A2 => p(0), A3 => p(1), A4 => p(2), Z => net_15);
	U58 : AND3 port map (A1 => g(0), A2 => p(1), A3 => p(2), Z => net_16);
	U59 : AND2 port map (A1 => g(1), A2 => p(2), Z => net_17);
	U60 : OR4 port map (A1 => net_15, A2 => net_16, A3 => net_17, A4 => g(2), Z => carry(3));
	U61 : AND3 port map (A1 => carry(0), A2 => p(0), A3 => p(1), Z => net_18);
	U62 : AND2 port map (A1 => g(0), A2 => p(1), Z => net_19);
	U63 : OR3 port map (A1 => net_18, A2 => net_19, A3 => g(1), Z => carry(2));
	U64 : AND2 port map (A1 => carry(0), A2 => p(0), Z => net_20);
	U65 : OR2 port map (A1 => net_20, A2 => g(0), Z => carry(1));
	carry(4) <= carry2(1);
	U66 : AND4 port map (A1 => carry(4), A2 => p(4), A3 => p(5), A4 => p(6), Z => net_21);
	U67 : AND3 port map (A1 => g(4), A2 => p(5), A3 => p(6), Z => net_22);
	U68 : AND2 port map (A1 => g(5), A2 => p(6), Z => net_23);
	U69 : OR4 port map (A1 => net_21, A2 => net_22, A3 => net_23, A4 => g(6), Z => carry(7));
	U70 : AND3 port map (A1 => carry(4), A2 => p(4), A3 => p(5), Z => net_24);
	U71 : AND2 port map (A1 => g(4), A2 => p(5), Z => net_25);
	U72 : OR3 port map (A1 => net_24, A2 => net_25, A3 => g(5), Z => carry(6));
	U73 : AND2 port map (A1 => carry(4), A2 => p(4), Z => net_26);
	U74 : OR2 port map (A1 => net_26, A2 => g(4), Z => carry(5));
	carry(8) <= carry2(2);
	U75 : AND4 port map (A1 => carry(8), A2 => p(8), A3 => p(9), A4 => p(10), Z => net_27);
	U76 : AND3 port map (A1 => g(8), A2 => p(9), A3 => p(10), Z => net_28);
	U77 : AND2 port map (A1 => g(9), A2 => p(10), Z => net_29);
	U78 : OR4 port map (A1 => net_27, A2 => net_28, A3 => net_29, A4 => g(10), Z => carry(11));
	U79 : AND3 port map (A1 => carry(8), A2 => p(8), A3 => p(9), Z => net_30);
	U80 : AND2 port map (A1 => g(8), A2 => p(9), Z => net_31);
	U81 : OR3 port map (A1 => net_30, A2 => net_31, A3 => g(9), Z => carry(10));
	U82 : AND2 port map (A1 => carry(8), A2 => p(8), Z => net_32);
	U83 : OR2 port map (A1 => net_32, A2 => g(8), Z => carry(9));
	carry(12) <= carry2(3);
	U84 : AND4 port map (A1 => carry(12), A2 => p(12), A3 => p(13), A4 => p(14), Z => net_33);
	U85 : AND3 port map (A1 => g(12), A2 => p(13), A3 => p(14), Z => net_34);
	U86 : AND2 port map (A1 => g(13), A2 => p(14), Z => net_35);
	U87 : OR4 port map (A1 => net_33, A2 => net_34, A3 => net_35, A4 => g(14), Z => carry(15));
	U88 : AND3 port map (A1 => carry(12), A2 => p(12), A3 => p(13), Z => net_36);
	U89 : AND2 port map (A1 => g(12), A2 => p(13), Z => net_37);
	U90 : OR3 port map (A1 => net_36, A2 => net_37, A3 => g(13), Z => carry(14));
	U91 : AND2 port map (A1 => carry(12), A2 => p(12), Z => net_38);
	U92 : OR2 port map (A1 => net_38, A2 => g(12), Z => carry(13));
	U93 : XOR2 port map (A1 => carry(0), A2 => p(0), Z => sum(0));
	U94 : XOR2 port map (A1 => carry(1), A2 => p(1), Z => sum(1));
	U95 : XOR2 port map (A1 => carry(2), A2 => p(2), Z => sum(2));
	U96 : XOR2 port map (A1 => carry(3), A2 => p(3), Z => sum(3));
	U97 : XOR2 port map (A1 => carry(4), A2 => p(4), Z => sum(4));
	U98 : XOR2 port map (A1 => carry(5), A2 => p(5), Z => sum(5));
	U99 : XOR2 port map (A1 => carry(6), A2 => p(6), Z => sum(6));
	U100 : XOR2 port map (A1 => carry(7), A2 => p(7), Z => sum(7));
	U101 : XOR2 port map (A1 => carry(8), A2 => p(8), Z => sum(8));
	U102 : XOR2 port map (A1 => carry(9), A2 => p(9), Z => sum(9));
	U103 : XOR2 port map (A1 => carry(10), A2 => p(10), Z => sum(10));
	U104 : XOR2 port map (A1 => carry(11), A2 => p(11), Z => sum(11));
	U105 : XOR2 port map (A1 => carry(12), A2 => p(12), Z => sum(12));
	U106 : XOR2 port map (A1 => carry(13), A2 => p(13), Z => sum(13));
	U107 : XOR2 port map (A1 => carry(14), A2 => p(14), Z => sum(14));
	U108 : XOR2 port map (A1 => carry(15), A2 => p(15), Z => sum(15));
end struct;
----------------------------------------------------------------------
