----------------------------------------------------------------------
entity adder64 is
	port (
		a        : in  std_logic_vector(63 downto 0);
		b        : in  std_logic_vector(63 downto 0);
		c_in     : in  std_logic;
		sum      : out std_logic_vector(63 downto 0)
	);
end adder64;
----------------------------------------------------------------------

----------------------------------------------------------------------
architecture struct of adder64 is
	signal p          : std_logic_vector(63 downto 0);
	signal g          : std_logic_vector(63 downto 0);
	signal carry      : std_logic_vector(63 downto 0);
	signal p2         : std_logic_vector(14 downto 0);
	signal g2         : std_logic_vector(14 downto 0);
	signal carry2     : std_logic_vector(15 downto 0);
	signal p3         : std_logic_vector(2 downto 0);
	signal g3         : std_logic_vector(2 downto 0);
	signal carry3     : std_logic_vector(3 downto 0);
	signal net_0      : std_logic;
	signal net_1      : std_logic;
	signal net_2      : std_logic;
	signal net_3      : std_logic;
	signal net_4      : std_logic;
	signal net_5      : std_logic;
	signal net_6      : std_logic;
	signal net_7      : std_logic;
	signal net_8      : std_logic;
	signal net_9      : std_logic;
	signal net_10     : std_logic;
	signal net_11     : std_logic;
	signal net_12     : std_logic;
	signal net_13     : std_logic;
	signal net_14     : std_logic;
	signal net_15     : std_logic;
	signal net_16     : std_logic;
	signal net_17     : std_logic;
	signal net_18     : std_logic;
	signal net_19     : std_logic;
	signal net_20     : std_logic;
	signal net_21     : std_logic;
	signal net_22     : std_logic;
	signal net_23     : std_logic;
	signal net_24     : std_logic;
	signal net_25     : std_logic;
	signal net_26     : std_logic;
	signal net_27     : std_logic;
	signal net_28     : std_logic;
	signal net_29     : std_logic;
	signal net_30     : std_logic;
	signal net_31     : std_logic;
	signal net_32     : std_logic;
	signal net_33     : std_logic;
	signal net_34     : std_logic;
	signal net_35     : std_logic;
	signal net_36     : std_logic;
	signal net_37     : std_logic;
	signal net_38     : std_logic;
	signal net_39     : std_logic;
	signal net_40     : std_logic;
	signal net_41     : std_logic;
	signal net_42     : std_logic;
	signal net_43     : std_logic;
	signal net_44     : std_logic;
	signal net_45     : std_logic;
	signal net_46     : std_logic;
	signal net_47     : std_logic;
	signal net_48     : std_logic;
	signal net_49     : std_logic;
	signal net_50     : std_logic;
	signal net_51     : std_logic;
	signal net_52     : std_logic;
	signal net_53     : std_logic;
	signal net_54     : std_logic;
	signal net_55     : std_logic;
	signal net_56     : std_logic;
	signal net_57     : std_logic;
	signal net_58     : std_logic;
	signal net_59     : std_logic;
	signal net_60     : std_logic;
	signal net_61     : std_logic;
	signal net_62     : std_logic;
	signal net_63     : std_logic;
	signal net_64     : std_logic;
	signal net_65     : std_logic;
	signal net_66     : std_logic;
	signal net_67     : std_logic;
	signal net_68     : std_logic;
	signal net_69     : std_logic;
	signal net_70     : std_logic;
	signal net_71     : std_logic;
	signal net_72     : std_logic;
	signal net_73     : std_logic;
	signal net_74     : std_logic;
	signal net_75     : std_logic;
	signal net_76     : std_logic;
	signal net_77     : std_logic;
	signal net_78     : std_logic;
	signal net_79     : std_logic;
	signal net_80     : std_logic;
	signal net_81     : std_logic;
	signal net_82     : std_logic;
	signal net_83     : std_logic;
	signal net_84     : std_logic;
	signal net_85     : std_logic;
	signal net_86     : std_logic;
	signal net_87     : std_logic;
	signal net_88     : std_logic;
	signal net_89     : std_logic;
	signal net_90     : std_logic;
	signal net_91     : std_logic;
	signal net_92     : std_logic;
	signal net_93     : std_logic;
	signal net_94     : std_logic;
	signal net_95     : std_logic;
	signal net_96     : std_logic;
	signal net_97     : std_logic;
	signal net_98     : std_logic;
	signal net_99     : std_logic;
	signal net_100    : std_logic;
	signal net_101    : std_logic;
	signal net_102    : std_logic;
	signal net_103    : std_logic;
	signal net_104    : std_logic;
	signal net_105    : std_logic;
	signal net_106    : std_logic;
	signal net_107    : std_logic;
	signal net_108    : std_logic;
	signal net_109    : std_logic;
	signal net_110    : std_logic;
	signal net_111    : std_logic;
	signal net_112    : std_logic;
	signal net_113    : std_logic;
	signal net_114    : std_logic;
	signal net_115    : std_logic;
	signal net_116    : std_logic;
	signal net_117    : std_logic;
	signal net_118    : std_logic;
	signal net_119    : std_logic;
	signal net_120    : std_logic;
	signal net_121    : std_logic;
	signal net_122    : std_logic;
	signal net_123    : std_logic;
	signal net_124    : std_logic;
	signal net_125    : std_logic;
	signal net_126    : std_logic;
	signal net_127    : std_logic;
	signal net_128    : std_logic;
	signal net_129    : std_logic;
	signal net_130    : std_logic;
	signal net_131    : std_logic;
	signal net_132    : std_logic;
	signal net_133    : std_logic;
	signal net_134    : std_logic;
	signal net_135    : std_logic;
	signal net_136    : std_logic;
	signal net_137    : std_logic;
	signal net_138    : std_logic;
	signal net_139    : std_logic;
	signal net_140    : std_logic;
	signal net_141    : std_logic;
	signal net_142    : std_logic;
	signal net_143    : std_logic;
	signal net_144    : std_logic;
	signal net_145    : std_logic;
	signal net_146    : std_logic;
	signal net_147    : std_logic;
	signal net_148    : std_logic;
	signal net_149    : std_logic;
	signal net_150    : std_logic;
	signal net_151    : std_logic;
	signal net_152    : std_logic;
	signal net_153    : std_logic;
	signal net_154    : std_logic;
	signal net_155    : std_logic;
	signal net_156    : std_logic;
	signal net_157    : std_logic;
	signal net_158    : std_logic;
	signal net_159    : std_logic;
	signal net_160    : std_logic;
	signal net_161    : std_logic;
	signal net_162    : std_logic;
	signal net_163    : std_logic;
	signal net_164    : std_logic;
	signal net_165    : std_logic;
	signal net_166    : std_logic;
	signal net_167    : std_logic;
	signal net_168    : std_logic;
	signal net_169    : std_logic;
	signal net_170    : std_logic;
	signal net_171    : std_logic;
	signal net_172    : std_logic;
	signal net_173    : std_logic;
	signal net_174    : std_logic;
	signal net_175    : std_logic;
	signal net_176    : std_logic;
	signal net_177    : std_logic;
	signal net_178    : std_logic;
	signal net_179    : std_logic;
begin
	carry(0) <= c_in;
	carry3(0) <= carry(0);
	carry2(0) <= carry3(0);
	carry2(4) <= carry3(1);
	carry2(8) <= carry3(2);
	carry2(12) <= carry3(3);
	carry(4) <= carry2(1);
	carry(8) <= carry2(2);
	carry(12) <= carry2(3);
	carry(16) <= carry2(4);
	carry(20) <= carry2(5);
	carry(24) <= carry2(6);
	carry(28) <= carry2(7);
	carry(32) <= carry2(8);
	carry(36) <= carry2(9);
	carry(40) <= carry2(10);
	carry(44) <= carry2(11);
	carry(48) <= carry2(12);
	carry(52) <= carry2(13);
	carry(56) <= carry2(14);
	carry(60) <= carry2(15);
	U1 : XOR2 port map(A1 => a(0), A2 => b(0), Z => p(0));
	U2 : AND2 port map(A1 => a(0), A2 => b(0), Z => g(0));
	U3 : XOR2 port map(A1 => a(1), A2 => b(1), Z => p(1));
	U4 : AND2 port map(A1 => a(1), A2 => b(1), Z => g(1));
	U5 : XOR2 port map(A1 => a(2), A2 => b(2), Z => p(2));
	U6 : AND2 port map(A1 => a(2), A2 => b(2), Z => g(2));
	U7 : XOR2 port map(A1 => a(3), A2 => b(3), Z => p(3));
	U8 : AND2 port map(A1 => a(3), A2 => b(3), Z => g(3));
	U9 : XOR2 port map(A1 => a(4), A2 => b(4), Z => p(4));
	U10 : AND2 port map(A1 => a(4), A2 => b(4), Z => g(4));
	U11 : XOR2 port map(A1 => a(5), A2 => b(5), Z => p(5));
	U12 : AND2 port map(A1 => a(5), A2 => b(5), Z => g(5));
	U13 : XOR2 port map(A1 => a(6), A2 => b(6), Z => p(6));
	U14 : AND2 port map(A1 => a(6), A2 => b(6), Z => g(6));
	U15 : XOR2 port map(A1 => a(7), A2 => b(7), Z => p(7));
	U16 : AND2 port map(A1 => a(7), A2 => b(7), Z => g(7));
	U17 : XOR2 port map(A1 => a(8), A2 => b(8), Z => p(8));
	U18 : AND2 port map(A1 => a(8), A2 => b(8), Z => g(8));
	U19 : XOR2 port map(A1 => a(9), A2 => b(9), Z => p(9));
	U20 : AND2 port map(A1 => a(9), A2 => b(9), Z => g(9));
	U21 : XOR2 port map(A1 => a(10), A2 => b(10), Z => p(10));
	U22 : AND2 port map(A1 => a(10), A2 => b(10), Z => g(10));
	U23 : XOR2 port map(A1 => a(11), A2 => b(11), Z => p(11));
	U24 : AND2 port map(A1 => a(11), A2 => b(11), Z => g(11));
	U25 : XOR2 port map(A1 => a(12), A2 => b(12), Z => p(12));
	U26 : AND2 port map(A1 => a(12), A2 => b(12), Z => g(12));
	U27 : XOR2 port map(A1 => a(13), A2 => b(13), Z => p(13));
	U28 : AND2 port map(A1 => a(13), A2 => b(13), Z => g(13));
	U29 : XOR2 port map(A1 => a(14), A2 => b(14), Z => p(14));
	U30 : AND2 port map(A1 => a(14), A2 => b(14), Z => g(14));
	U31 : XOR2 port map(A1 => a(15), A2 => b(15), Z => p(15));
	U32 : AND2 port map(A1 => a(15), A2 => b(15), Z => g(15));
	U33 : XOR2 port map(A1 => a(16), A2 => b(16), Z => p(16));
	U34 : AND2 port map(A1 => a(16), A2 => b(16), Z => g(16));
	U35 : XOR2 port map(A1 => a(17), A2 => b(17), Z => p(17));
	U36 : AND2 port map(A1 => a(17), A2 => b(17), Z => g(17));
	U37 : XOR2 port map(A1 => a(18), A2 => b(18), Z => p(18));
	U38 : AND2 port map(A1 => a(18), A2 => b(18), Z => g(18));
	U39 : XOR2 port map(A1 => a(19), A2 => b(19), Z => p(19));
	U40 : AND2 port map(A1 => a(19), A2 => b(19), Z => g(19));
	U41 : XOR2 port map(A1 => a(20), A2 => b(20), Z => p(20));
	U42 : AND2 port map(A1 => a(20), A2 => b(20), Z => g(20));
	U43 : XOR2 port map(A1 => a(21), A2 => b(21), Z => p(21));
	U44 : AND2 port map(A1 => a(21), A2 => b(21), Z => g(21));
	U45 : XOR2 port map(A1 => a(22), A2 => b(22), Z => p(22));
	U46 : AND2 port map(A1 => a(22), A2 => b(22), Z => g(22));
	U47 : XOR2 port map(A1 => a(23), A2 => b(23), Z => p(23));
	U48 : AND2 port map(A1 => a(23), A2 => b(23), Z => g(23));
	U49 : XOR2 port map(A1 => a(24), A2 => b(24), Z => p(24));
	U50 : AND2 port map(A1 => a(24), A2 => b(24), Z => g(24));
	U51 : XOR2 port map(A1 => a(25), A2 => b(25), Z => p(25));
	U52 : AND2 port map(A1 => a(25), A2 => b(25), Z => g(25));
	U53 : XOR2 port map(A1 => a(26), A2 => b(26), Z => p(26));
	U54 : AND2 port map(A1 => a(26), A2 => b(26), Z => g(26));
	U55 : XOR2 port map(A1 => a(27), A2 => b(27), Z => p(27));
	U56 : AND2 port map(A1 => a(27), A2 => b(27), Z => g(27));
	U57 : XOR2 port map(A1 => a(28), A2 => b(28), Z => p(28));
	U58 : AND2 port map(A1 => a(28), A2 => b(28), Z => g(28));
	U59 : XOR2 port map(A1 => a(29), A2 => b(29), Z => p(29));
	U60 : AND2 port map(A1 => a(29), A2 => b(29), Z => g(29));
	U61 : XOR2 port map(A1 => a(30), A2 => b(30), Z => p(30));
	U62 : AND2 port map(A1 => a(30), A2 => b(30), Z => g(30));
	U63 : XOR2 port map(A1 => a(31), A2 => b(31), Z => p(31));
	U64 : AND2 port map(A1 => a(31), A2 => b(31), Z => g(31));
	U65 : XOR2 port map(A1 => a(32), A2 => b(32), Z => p(32));
	U66 : AND2 port map(A1 => a(32), A2 => b(32), Z => g(32));
	U67 : XOR2 port map(A1 => a(33), A2 => b(33), Z => p(33));
	U68 : AND2 port map(A1 => a(33), A2 => b(33), Z => g(33));
	U69 : XOR2 port map(A1 => a(34), A2 => b(34), Z => p(34));
	U70 : AND2 port map(A1 => a(34), A2 => b(34), Z => g(34));
	U71 : XOR2 port map(A1 => a(35), A2 => b(35), Z => p(35));
	U72 : AND2 port map(A1 => a(35), A2 => b(35), Z => g(35));
	U73 : XOR2 port map(A1 => a(36), A2 => b(36), Z => p(36));
	U74 : AND2 port map(A1 => a(36), A2 => b(36), Z => g(36));
	U75 : XOR2 port map(A1 => a(37), A2 => b(37), Z => p(37));
	U76 : AND2 port map(A1 => a(37), A2 => b(37), Z => g(37));
	U77 : XOR2 port map(A1 => a(38), A2 => b(38), Z => p(38));
	U78 : AND2 port map(A1 => a(38), A2 => b(38), Z => g(38));
	U79 : XOR2 port map(A1 => a(39), A2 => b(39), Z => p(39));
	U80 : AND2 port map(A1 => a(39), A2 => b(39), Z => g(39));
	U81 : XOR2 port map(A1 => a(40), A2 => b(40), Z => p(40));
	U82 : AND2 port map(A1 => a(40), A2 => b(40), Z => g(40));
	U83 : XOR2 port map(A1 => a(41), A2 => b(41), Z => p(41));
	U84 : AND2 port map(A1 => a(41), A2 => b(41), Z => g(41));
	U85 : XOR2 port map(A1 => a(42), A2 => b(42), Z => p(42));
	U86 : AND2 port map(A1 => a(42), A2 => b(42), Z => g(42));
	U87 : XOR2 port map(A1 => a(43), A2 => b(43), Z => p(43));
	U88 : AND2 port map(A1 => a(43), A2 => b(43), Z => g(43));
	U89 : XOR2 port map(A1 => a(44), A2 => b(44), Z => p(44));
	U90 : AND2 port map(A1 => a(44), A2 => b(44), Z => g(44));
	U91 : XOR2 port map(A1 => a(45), A2 => b(45), Z => p(45));
	U92 : AND2 port map(A1 => a(45), A2 => b(45), Z => g(45));
	U93 : XOR2 port map(A1 => a(46), A2 => b(46), Z => p(46));
	U94 : AND2 port map(A1 => a(46), A2 => b(46), Z => g(46));
	U95 : XOR2 port map(A1 => a(47), A2 => b(47), Z => p(47));
	U96 : AND2 port map(A1 => a(47), A2 => b(47), Z => g(47));
	U97 : XOR2 port map(A1 => a(48), A2 => b(48), Z => p(48));
	U98 : AND2 port map(A1 => a(48), A2 => b(48), Z => g(48));
	U99 : XOR2 port map(A1 => a(49), A2 => b(49), Z => p(49));
	U100 : AND2 port map(A1 => a(49), A2 => b(49), Z => g(49));
	U101 : XOR2 port map(A1 => a(50), A2 => b(50), Z => p(50));
	U102 : AND2 port map(A1 => a(50), A2 => b(50), Z => g(50));
	U103 : XOR2 port map(A1 => a(51), A2 => b(51), Z => p(51));
	U104 : AND2 port map(A1 => a(51), A2 => b(51), Z => g(51));
	U105 : XOR2 port map(A1 => a(52), A2 => b(52), Z => p(52));
	U106 : AND2 port map(A1 => a(52), A2 => b(52), Z => g(52));
	U107 : XOR2 port map(A1 => a(53), A2 => b(53), Z => p(53));
	U108 : AND2 port map(A1 => a(53), A2 => b(53), Z => g(53));
	U109 : XOR2 port map(A1 => a(54), A2 => b(54), Z => p(54));
	U110 : AND2 port map(A1 => a(54), A2 => b(54), Z => g(54));
	U111 : XOR2 port map(A1 => a(55), A2 => b(55), Z => p(55));
	U112 : AND2 port map(A1 => a(55), A2 => b(55), Z => g(55));
	U113 : XOR2 port map(A1 => a(56), A2 => b(56), Z => p(56));
	U114 : AND2 port map(A1 => a(56), A2 => b(56), Z => g(56));
	U115 : XOR2 port map(A1 => a(57), A2 => b(57), Z => p(57));
	U116 : AND2 port map(A1 => a(57), A2 => b(57), Z => g(57));
	U117 : XOR2 port map(A1 => a(58), A2 => b(58), Z => p(58));
	U118 : AND2 port map(A1 => a(58), A2 => b(58), Z => g(58));
	U119 : XOR2 port map(A1 => a(59), A2 => b(59), Z => p(59));
	U120 : AND2 port map(A1 => a(59), A2 => b(59), Z => g(59));
	U121 : XOR2 port map(A1 => a(60), A2 => b(60), Z => p(60));
	U122 : AND2 port map(A1 => a(60), A2 => b(60), Z => g(60));
	U123 : XOR2 port map(A1 => a(61), A2 => b(61), Z => p(61));
	U124 : AND2 port map(A1 => a(61), A2 => b(61), Z => g(61));
	U125 : XOR2 port map(A1 => a(62), A2 => b(62), Z => p(62));
	U126 : AND2 port map(A1 => a(62), A2 => b(62), Z => g(62));
	U127 : XOR2 port map(A1 => a(63), A2 => b(63), Z => p(63));
	U128 : AND2 port map(A1 => a(63), A2 => b(63), Z => g(63));
	U129 : AND4 port map(A1 => p(0), A2 => p(1), A3 => p(2), A4 => p(3), Z => p2(0));
	U130 : AND4 port map(A1 => p(4), A2 => p(5), A3 => p(6), A4 => p(7), Z => p2(1));
	U131 : AND4 port map(A1 => p(8), A2 => p(9), A3 => p(10), A4 => p(11), Z => p2(2));
	U132 : AND4 port map(A1 => p(12), A2 => p(13), A3 => p(14), A4 => p(15), Z => p2(3));
	U133 : AND4 port map(A1 => p(16), A2 => p(17), A3 => p(18), A4 => p(19), Z => p2(4));
	U134 : AND4 port map(A1 => p(20), A2 => p(21), A3 => p(22), A4 => p(23), Z => p2(5));
	U135 : AND4 port map(A1 => p(24), A2 => p(25), A3 => p(26), A4 => p(27), Z => p2(6));
	U136 : AND4 port map(A1 => p(28), A2 => p(29), A3 => p(30), A4 => p(31), Z => p2(7));
	U137 : AND4 port map(A1 => p(32), A2 => p(33), A3 => p(34), A4 => p(35), Z => p2(8));
	U138 : AND4 port map(A1 => p(36), A2 => p(37), A3 => p(38), A4 => p(39), Z => p2(9));
	U139 : AND4 port map(A1 => p(40), A2 => p(41), A3 => p(42), A4 => p(43), Z => p2(10));
	U140 : AND4 port map(A1 => p(44), A2 => p(45), A3 => p(46), A4 => p(47), Z => p2(11));
	U141 : AND4 port map(A1 => p(48), A2 => p(49), A3 => p(50), A4 => p(51), Z => p2(12));
	U142 : AND4 port map(A1 => p(52), A2 => p(53), A3 => p(54), A4 => p(55), Z => p2(13));
	U143 : AND4 port map(A1 => p(56), A2 => p(57), A3 => p(58), A4 => p(59), Z => p2(14));
	U144 : AND4 port map(A1 => g(0), A2 => p(1), A3 => p(2), A4 => p(3), Z => net_0);
	U145 : AND3 port map(A1 => g(1), A2 => p(2), A3 => p(3), Z => net_1);
	U146 : AND2 port map(A1 => g(2), A2 => p(3), Z => net_2);
	U147 : OR4 port map(A1 => net_0, A2 => net_1, A3 => net_2, A4 => g(3), Z => g2(0));
	U148 : AND4 port map(A1 => g(4), A2 => p(5), A3 => p(6), A4 => p(7), Z => net_3);
	U149 : AND3 port map(A1 => g(5), A2 => p(6), A3 => p(7), Z => net_4);
	U150 : AND2 port map(A1 => g(6), A2 => p(7), Z => net_5);
	U151 : OR4 port map(A1 => net_3, A2 => net_4, A3 => net_5, A4 => g(7), Z => g2(1));
	U152 : AND4 port map(A1 => g(8), A2 => p(9), A3 => p(10), A4 => p(11), Z => net_6);
	U153 : AND3 port map(A1 => g(9), A2 => p(10), A3 => p(11), Z => net_7);
	U154 : AND2 port map(A1 => g(10), A2 => p(11), Z => net_8);
	U155 : OR4 port map(A1 => net_6, A2 => net_7, A3 => net_8, A4 => g(11), Z => g2(2));
	U156 : AND4 port map(A1 => g(12), A2 => p(13), A3 => p(14), A4 => p(15), Z => net_9);
	U157 : AND3 port map(A1 => g(13), A2 => p(14), A3 => p(15), Z => net_10);
	U158 : AND2 port map(A1 => g(14), A2 => p(15), Z => net_11);
	U159 : OR4 port map(A1 => net_9, A2 => net_10, A3 => net_11, A4 => g(15), Z => g2(3));
	U160 : AND4 port map(A1 => g(16), A2 => p(17), A3 => p(18), A4 => p(19), Z => net_12);
	U161 : AND3 port map(A1 => g(17), A2 => p(18), A3 => p(19), Z => net_13);
	U162 : AND2 port map(A1 => g(18), A2 => p(19), Z => net_14);
	U163 : OR4 port map(A1 => net_12, A2 => net_13, A3 => net_14, A4 => g(19), Z => g2(4));
	U164 : AND4 port map(A1 => g(20), A2 => p(21), A3 => p(22), A4 => p(23), Z => net_15);
	U165 : AND3 port map(A1 => g(21), A2 => p(22), A3 => p(23), Z => net_16);
	U166 : AND2 port map(A1 => g(22), A2 => p(23), Z => net_17);
	U167 : OR4 port map(A1 => net_15, A2 => net_16, A3 => net_17, A4 => g(23), Z => g2(5));
	U168 : AND4 port map(A1 => g(24), A2 => p(25), A3 => p(26), A4 => p(27), Z => net_18);
	U169 : AND3 port map(A1 => g(25), A2 => p(26), A3 => p(27), Z => net_19);
	U170 : AND2 port map(A1 => g(26), A2 => p(27), Z => net_20);
	U171 : OR4 port map(A1 => net_18, A2 => net_19, A3 => net_20, A4 => g(27), Z => g2(6));
	U172 : AND4 port map(A1 => g(28), A2 => p(29), A3 => p(30), A4 => p(31), Z => net_21);
	U173 : AND3 port map(A1 => g(29), A2 => p(30), A3 => p(31), Z => net_22);
	U174 : AND2 port map(A1 => g(30), A2 => p(31), Z => net_23);
	U175 : OR4 port map(A1 => net_21, A2 => net_22, A3 => net_23, A4 => g(31), Z => g2(7));
	U176 : AND4 port map(A1 => g(32), A2 => p(33), A3 => p(34), A4 => p(35), Z => net_24);
	U177 : AND3 port map(A1 => g(33), A2 => p(34), A3 => p(35), Z => net_25);
	U178 : AND2 port map(A1 => g(34), A2 => p(35), Z => net_26);
	U179 : OR4 port map(A1 => net_24, A2 => net_25, A3 => net_26, A4 => g(35), Z => g2(8));
	U180 : AND4 port map(A1 => g(36), A2 => p(37), A3 => p(38), A4 => p(39), Z => net_27);
	U181 : AND3 port map(A1 => g(37), A2 => p(38), A3 => p(39), Z => net_28);
	U182 : AND2 port map(A1 => g(38), A2 => p(39), Z => net_29);
	U183 : OR4 port map(A1 => net_27, A2 => net_28, A3 => net_29, A4 => g(39), Z => g2(9));
	U184 : AND4 port map(A1 => g(40), A2 => p(41), A3 => p(42), A4 => p(43), Z => net_30);
	U185 : AND3 port map(A1 => g(41), A2 => p(42), A3 => p(43), Z => net_31);
	U186 : AND2 port map(A1 => g(42), A2 => p(43), Z => net_32);
	U187 : OR4 port map(A1 => net_30, A2 => net_31, A3 => net_32, A4 => g(43), Z => g2(10));
	U188 : AND4 port map(A1 => g(44), A2 => p(45), A3 => p(46), A4 => p(47), Z => net_33);
	U189 : AND3 port map(A1 => g(45), A2 => p(46), A3 => p(47), Z => net_34);
	U190 : AND2 port map(A1 => g(46), A2 => p(47), Z => net_35);
	U191 : OR4 port map(A1 => net_33, A2 => net_34, A3 => net_35, A4 => g(47), Z => g2(11));
	U192 : AND4 port map(A1 => g(48), A2 => p(49), A3 => p(50), A4 => p(51), Z => net_36);
	U193 : AND3 port map(A1 => g(49), A2 => p(50), A3 => p(51), Z => net_37);
	U194 : AND2 port map(A1 => g(50), A2 => p(51), Z => net_38);
	U195 : OR4 port map(A1 => net_36, A2 => net_37, A3 => net_38, A4 => g(51), Z => g2(12));
	U196 : AND4 port map(A1 => g(52), A2 => p(53), A3 => p(54), A4 => p(55), Z => net_39);
	U197 : AND3 port map(A1 => g(53), A2 => p(54), A3 => p(55), Z => net_40);
	U198 : AND2 port map(A1 => g(54), A2 => p(55), Z => net_41);
	U199 : OR4 port map(A1 => net_39, A2 => net_40, A3 => net_41, A4 => g(55), Z => g2(13));
	U200 : AND4 port map(A1 => g(56), A2 => p(57), A3 => p(58), A4 => p(59), Z => net_42);
	U201 : AND3 port map(A1 => g(57), A2 => p(58), A3 => p(59), Z => net_43);
	U202 : AND2 port map(A1 => g(58), A2 => p(59), Z => net_44);
	U203 : OR4 port map(A1 => net_42, A2 => net_43, A3 => net_44, A4 => g(59), Z => g2(14));
	U204 : AND4 port map(A1 => p2(0), A2 => p2(1), A3 => p2(2), A4 => p2(3), Z => p3(0));
	U205 : AND4 port map(A1 => p2(4), A2 => p2(5), A3 => p2(6), A4 => p2(7), Z => p3(1));
	U206 : AND4 port map(A1 => p2(8), A2 => p2(9), A3 => p2(10), A4 => p2(11), Z => p3(2));
	U207 : AND4 port map(A1 => g2(0), A2 => p2(1), A3 => p2(2), A4 => p2(3), Z => net_45);
	U208 : AND3 port map(A1 => g2(1), A2 => p2(2), A3 => p2(3), Z => net_46);
	U209 : AND2 port map(A1 => g2(2), A2 => p2(3), Z => net_47);
	U210 : OR4 port map(A1 => net_45, A2 => net_46, A3 => net_47, A4 => g2(3), Z => g3(0));
	U211 : AND4 port map(A1 => g2(4), A2 => p2(5), A3 => p2(6), A4 => p2(7), Z => net_48);
	U212 : AND3 port map(A1 => g2(5), A2 => p2(6), A3 => p2(7), Z => net_49);
	U213 : AND2 port map(A1 => g2(6), A2 => p2(7), Z => net_50);
	U214 : OR4 port map(A1 => net_48, A2 => net_49, A3 => net_50, A4 => g2(7), Z => g3(1));
	U215 : AND4 port map(A1 => g2(8), A2 => p2(9), A3 => p2(10), A4 => p2(11), Z => net_51);
	U216 : AND3 port map(A1 => g2(9), A2 => p2(10), A3 => p2(11), Z => net_52);
	U217 : AND2 port map(A1 => g2(10), A2 => p2(11), Z => net_53);
	U218 : OR4 port map(A1 => net_51, A2 => net_52, A3 => net_53, A4 => g2(11), Z => g3(2));
	U219 : AND4 port map(A1 => carry3(0), A2 => p3(0), A3 => p3(1), A4 => p3(2), Z => net_54);
	U220 : AND3 port map(A1 => g3(0), A2 => p3(1), A3 => p3(2), Z => net_55);
	U221 : AND2 port map(A1 => g3(1), A2 => p3(2), Z => net_56);
	U222 : OR4 port map(A1 => net_54, A2 => net_55, A3 => net_56, A4 => g3(2), Z => carry3(3));
	U223 : AND3 port map(A1 => carry3(0), A2 => p3(0), A3 => p3(1), Z => net_57);
	U224 : AND2 port map(A1 => g3(0), A2 => p3(1), Z => net_58);
	U225 : OR3 port map(A1 => net_57, A2 => net_58, A3 => g3(1), Z => carry3(2));
	U226 : AND2 port map(A1 => carry3(0), A2 => p3(0), Z => net_59);
	U227 : OR2 port map(A1 => net_59, A2 => g3(0), Z => carry3(1));
	U228 : AND4 port map(A1 => carry2(0), A2 => p2(0), A3 => p2(1), A4 => p2(2), Z => net_60);
	U229 : AND3 port map(A1 => g2(0), A2 => p2(1), A3 => p2(2), Z => net_61);
	U230 : AND2 port map(A1 => g2(1), A2 => p2(2), Z => net_62);
	U231 : OR4 port map(A1 => net_60, A2 => net_61, A3 => net_62, A4 => g2(2), Z => carry2(3));
	U232 : AND3 port map(A1 => carry2(0), A2 => p2(0), A3 => p2(1), Z => net_63);
	U233 : AND2 port map(A1 => g2(0), A2 => p2(1), Z => net_64);
	U234 : OR3 port map(A1 => net_63, A2 => net_64, A3 => g2(1), Z => carry2(2));
	U235 : AND2 port map(A1 => carry2(0), A2 => p2(0), Z => net_65);
	U236 : OR2 port map(A1 => net_65, A2 => g2(0), Z => carry2(1));
	U237 : AND4 port map(A1 => carry2(4), A2 => p2(4), A3 => p2(5), A4 => p2(6), Z => net_66);
	U238 : AND3 port map(A1 => g2(4), A2 => p2(5), A3 => p2(6), Z => net_67);
	U239 : AND2 port map(A1 => g2(5), A2 => p2(6), Z => net_68);
	U240 : OR4 port map(A1 => net_66, A2 => net_67, A3 => net_68, A4 => g2(6), Z => carry2(7));
	U241 : AND3 port map(A1 => carry2(4), A2 => p2(4), A3 => p2(5), Z => net_69);
	U242 : AND2 port map(A1 => g2(4), A2 => p2(5), Z => net_70);
	U243 : OR3 port map(A1 => net_69, A2 => net_70, A3 => g2(5), Z => carry2(6));
	U244 : AND2 port map(A1 => carry2(4), A2 => p2(4), Z => net_71);
	U245 : OR2 port map(A1 => net_71, A2 => g2(4), Z => carry2(5));
	U246 : AND4 port map(A1 => carry2(8), A2 => p2(8), A3 => p2(9), A4 => p2(10), Z => net_72);
	U247 : AND3 port map(A1 => g2(8), A2 => p2(9), A3 => p2(10), Z => net_73);
	U248 : AND2 port map(A1 => g2(9), A2 => p2(10), Z => net_74);
	U249 : OR4 port map(A1 => net_72, A2 => net_73, A3 => net_74, A4 => g2(10), Z => carry2(11));
	U250 : AND3 port map(A1 => carry2(8), A2 => p2(8), A3 => p2(9), Z => net_75);
	U251 : AND2 port map(A1 => g2(8), A2 => p2(9), Z => net_76);
	U252 : OR3 port map(A1 => net_75, A2 => net_76, A3 => g2(9), Z => carry2(10));
	U253 : AND2 port map(A1 => carry2(8), A2 => p2(8), Z => net_77);
	U254 : OR2 port map(A1 => net_77, A2 => g2(8), Z => carry2(9));
	U255 : AND4 port map(A1 => carry2(12), A2 => p2(12), A3 => p2(13), A4 => p2(14), Z => net_78);
	U256 : AND3 port map(A1 => g2(12), A2 => p2(13), A3 => p2(14), Z => net_79);
	U257 : AND2 port map(A1 => g2(13), A2 => p2(14), Z => net_80);
	U258 : OR4 port map(A1 => net_78, A2 => net_79, A3 => net_80, A4 => g2(14), Z => carry2(15));
	U259 : AND3 port map(A1 => carry2(12), A2 => p2(12), A3 => p2(13), Z => net_81);
	U260 : AND2 port map(A1 => g2(12), A2 => p2(13), Z => net_82);
	U261 : OR3 port map(A1 => net_81, A2 => net_82, A3 => g2(13), Z => carry2(14));
	U262 : AND2 port map(A1 => carry2(12), A2 => p2(12), Z => net_83);
	U263 : OR2 port map(A1 => net_83, A2 => g2(12), Z => carry2(13));
	U264 : AND4 port map(A1 => carry(0), A2 => p(0), A3 => p(1), A4 => p(2), Z => net_84);
	U265 : AND3 port map(A1 => g(0), A2 => p(1), A3 => p(2), Z => net_85);
	U266 : AND2 port map(A1 => g(1), A2 => p(2), Z => net_86);
	U267 : OR4 port map(A1 => net_84, A2 => net_85, A3 => net_86, A4 => g(2), Z => carry(3));
	U268 : AND3 port map(A1 => carry(0), A2 => p(0), A3 => p(1), Z => net_87);
	U269 : AND2 port map(A1 => g(0), A2 => p(1), Z => net_88);
	U270 : OR3 port map(A1 => net_87, A2 => net_88, A3 => g(1), Z => carry(2));
	U271 : AND2 port map(A1 => carry(0), A2 => p(0), Z => net_89);
	U272 : OR2 port map(A1 => net_89, A2 => g(0), Z => carry(1));
	U273 : AND4 port map(A1 => carry(4), A2 => p(4), A3 => p(5), A4 => p(6), Z => net_90);
	U274 : AND3 port map(A1 => g(4), A2 => p(5), A3 => p(6), Z => net_91);
	U275 : AND2 port map(A1 => g(5), A2 => p(6), Z => net_92);
	U276 : OR4 port map(A1 => net_90, A2 => net_91, A3 => net_92, A4 => g(6), Z => carry(7));
	U277 : AND3 port map(A1 => carry(4), A2 => p(4), A3 => p(5), Z => net_93);
	U278 : AND2 port map(A1 => g(4), A2 => p(5), Z => net_94);
	U279 : OR3 port map(A1 => net_93, A2 => net_94, A3 => g(5), Z => carry(6));
	U280 : AND2 port map(A1 => carry(4), A2 => p(4), Z => net_95);
	U281 : OR2 port map(A1 => net_95, A2 => g(4), Z => carry(5));
	U282 : AND4 port map(A1 => carry(8), A2 => p(8), A3 => p(9), A4 => p(10), Z => net_96);
	U283 : AND3 port map(A1 => g(8), A2 => p(9), A3 => p(10), Z => net_97);
	U284 : AND2 port map(A1 => g(9), A2 => p(10), Z => net_98);
	U285 : OR4 port map(A1 => net_96, A2 => net_97, A3 => net_98, A4 => g(10), Z => carry(11));
	U286 : AND3 port map(A1 => carry(8), A2 => p(8), A3 => p(9), Z => net_99);
	U287 : AND2 port map(A1 => g(8), A2 => p(9), Z => net_100);
	U288 : OR3 port map(A1 => net_99, A2 => net_100, A3 => g(9), Z => carry(10));
	U289 : AND2 port map(A1 => carry(8), A2 => p(8), Z => net_101);
	U290 : OR2 port map(A1 => net_101, A2 => g(8), Z => carry(9));
	U291 : AND4 port map(A1 => carry(12), A2 => p(12), A3 => p(13), A4 => p(14), Z => net_102);
	U292 : AND3 port map(A1 => g(12), A2 => p(13), A3 => p(14), Z => net_103);
	U293 : AND2 port map(A1 => g(13), A2 => p(14), Z => net_104);
	U294 : OR4 port map(A1 => net_102, A2 => net_103, A3 => net_104, A4 => g(14), Z => carry(15));
	U295 : AND3 port map(A1 => carry(12), A2 => p(12), A3 => p(13), Z => net_105);
	U296 : AND2 port map(A1 => g(12), A2 => p(13), Z => net_106);
	U297 : OR3 port map(A1 => net_105, A2 => net_106, A3 => g(13), Z => carry(14));
	U298 : AND2 port map(A1 => carry(12), A2 => p(12), Z => net_107);
	U299 : OR2 port map(A1 => net_107, A2 => g(12), Z => carry(13));
	U300 : AND4 port map(A1 => carry(16), A2 => p(16), A3 => p(17), A4 => p(18), Z => net_108);
	U301 : AND3 port map(A1 => g(16), A2 => p(17), A3 => p(18), Z => net_109);
	U302 : AND2 port map(A1 => g(17), A2 => p(18), Z => net_110);
	U303 : OR4 port map(A1 => net_108, A2 => net_109, A3 => net_110, A4 => g(18), Z => carry(19));
	U304 : AND3 port map(A1 => carry(16), A2 => p(16), A3 => p(17), Z => net_111);
	U305 : AND2 port map(A1 => g(16), A2 => p(17), Z => net_112);
	U306 : OR3 port map(A1 => net_111, A2 => net_112, A3 => g(17), Z => carry(18));
	U307 : AND2 port map(A1 => carry(16), A2 => p(16), Z => net_113);
	U308 : OR2 port map(A1 => net_113, A2 => g(16), Z => carry(17));
	U309 : AND4 port map(A1 => carry(20), A2 => p(20), A3 => p(21), A4 => p(22), Z => net_114);
	U310 : AND3 port map(A1 => g(20), A2 => p(21), A3 => p(22), Z => net_115);
	U311 : AND2 port map(A1 => g(21), A2 => p(22), Z => net_116);
	U312 : OR4 port map(A1 => net_114, A2 => net_115, A3 => net_116, A4 => g(22), Z => carry(23));
	U313 : AND3 port map(A1 => carry(20), A2 => p(20), A3 => p(21), Z => net_117);
	U314 : AND2 port map(A1 => g(20), A2 => p(21), Z => net_118);
	U315 : OR3 port map(A1 => net_117, A2 => net_118, A3 => g(21), Z => carry(22));
	U316 : AND2 port map(A1 => carry(20), A2 => p(20), Z => net_119);
	U317 : OR2 port map(A1 => net_119, A2 => g(20), Z => carry(21));
	U318 : AND4 port map(A1 => carry(24), A2 => p(24), A3 => p(25), A4 => p(26), Z => net_120);
	U319 : AND3 port map(A1 => g(24), A2 => p(25), A3 => p(26), Z => net_121);
	U320 : AND2 port map(A1 => g(25), A2 => p(26), Z => net_122);
	U321 : OR4 port map(A1 => net_120, A2 => net_121, A3 => net_122, A4 => g(26), Z => carry(27));
	U322 : AND3 port map(A1 => carry(24), A2 => p(24), A3 => p(25), Z => net_123);
	U323 : AND2 port map(A1 => g(24), A2 => p(25), Z => net_124);
	U324 : OR3 port map(A1 => net_123, A2 => net_124, A3 => g(25), Z => carry(26));
	U325 : AND2 port map(A1 => carry(24), A2 => p(24), Z => net_125);
	U326 : OR2 port map(A1 => net_125, A2 => g(24), Z => carry(25));
	U327 : AND4 port map(A1 => carry(28), A2 => p(28), A3 => p(29), A4 => p(30), Z => net_126);
	U328 : AND3 port map(A1 => g(28), A2 => p(29), A3 => p(30), Z => net_127);
	U329 : AND2 port map(A1 => g(29), A2 => p(30), Z => net_128);
	U330 : OR4 port map(A1 => net_126, A2 => net_127, A3 => net_128, A4 => g(30), Z => carry(31));
	U331 : AND3 port map(A1 => carry(28), A2 => p(28), A3 => p(29), Z => net_129);
	U332 : AND2 port map(A1 => g(28), A2 => p(29), Z => net_130);
	U333 : OR3 port map(A1 => net_129, A2 => net_130, A3 => g(29), Z => carry(30));
	U334 : AND2 port map(A1 => carry(28), A2 => p(28), Z => net_131);
	U335 : OR2 port map(A1 => net_131, A2 => g(28), Z => carry(29));
	U336 : AND4 port map(A1 => carry(32), A2 => p(32), A3 => p(33), A4 => p(34), Z => net_132);
	U337 : AND3 port map(A1 => g(32), A2 => p(33), A3 => p(34), Z => net_133);
	U338 : AND2 port map(A1 => g(33), A2 => p(34), Z => net_134);
	U339 : OR4 port map(A1 => net_132, A2 => net_133, A3 => net_134, A4 => g(34), Z => carry(35));
	U340 : AND3 port map(A1 => carry(32), A2 => p(32), A3 => p(33), Z => net_135);
	U341 : AND2 port map(A1 => g(32), A2 => p(33), Z => net_136);
	U342 : OR3 port map(A1 => net_135, A2 => net_136, A3 => g(33), Z => carry(34));
	U343 : AND2 port map(A1 => carry(32), A2 => p(32), Z => net_137);
	U344 : OR2 port map(A1 => net_137, A2 => g(32), Z => carry(33));
	U345 : AND4 port map(A1 => carry(36), A2 => p(36), A3 => p(37), A4 => p(38), Z => net_138);
	U346 : AND3 port map(A1 => g(36), A2 => p(37), A3 => p(38), Z => net_139);
	U347 : AND2 port map(A1 => g(37), A2 => p(38), Z => net_140);
	U348 : OR4 port map(A1 => net_138, A2 => net_139, A3 => net_140, A4 => g(38), Z => carry(39));
	U349 : AND3 port map(A1 => carry(36), A2 => p(36), A3 => p(37), Z => net_141);
	U350 : AND2 port map(A1 => g(36), A2 => p(37), Z => net_142);
	U351 : OR3 port map(A1 => net_141, A2 => net_142, A3 => g(37), Z => carry(38));
	U352 : AND2 port map(A1 => carry(36), A2 => p(36), Z => net_143);
	U353 : OR2 port map(A1 => net_143, A2 => g(36), Z => carry(37));
	U354 : AND4 port map(A1 => carry(40), A2 => p(40), A3 => p(41), A4 => p(42), Z => net_144);
	U355 : AND3 port map(A1 => g(40), A2 => p(41), A3 => p(42), Z => net_145);
	U356 : AND2 port map(A1 => g(41), A2 => p(42), Z => net_146);
	U357 : OR4 port map(A1 => net_144, A2 => net_145, A3 => net_146, A4 => g(42), Z => carry(43));
	U358 : AND3 port map(A1 => carry(40), A2 => p(40), A3 => p(41), Z => net_147);
	U359 : AND2 port map(A1 => g(40), A2 => p(41), Z => net_148);
	U360 : OR3 port map(A1 => net_147, A2 => net_148, A3 => g(41), Z => carry(42));
	U361 : AND2 port map(A1 => carry(40), A2 => p(40), Z => net_149);
	U362 : OR2 port map(A1 => net_149, A2 => g(40), Z => carry(41));
	U363 : AND4 port map(A1 => carry(44), A2 => p(44), A3 => p(45), A4 => p(46), Z => net_150);
	U364 : AND3 port map(A1 => g(44), A2 => p(45), A3 => p(46), Z => net_151);
	U365 : AND2 port map(A1 => g(45), A2 => p(46), Z => net_152);
	U366 : OR4 port map(A1 => net_150, A2 => net_151, A3 => net_152, A4 => g(46), Z => carry(47));
	U367 : AND3 port map(A1 => carry(44), A2 => p(44), A3 => p(45), Z => net_153);
	U368 : AND2 port map(A1 => g(44), A2 => p(45), Z => net_154);
	U369 : OR3 port map(A1 => net_153, A2 => net_154, A3 => g(45), Z => carry(46));
	U370 : AND2 port map(A1 => carry(44), A2 => p(44), Z => net_155);
	U371 : OR2 port map(A1 => net_155, A2 => g(44), Z => carry(45));
	U372 : AND4 port map(A1 => carry(48), A2 => p(48), A3 => p(49), A4 => p(50), Z => net_156);
	U373 : AND3 port map(A1 => g(48), A2 => p(49), A3 => p(50), Z => net_157);
	U374 : AND2 port map(A1 => g(49), A2 => p(50), Z => net_158);
	U375 : OR4 port map(A1 => net_156, A2 => net_157, A3 => net_158, A4 => g(50), Z => carry(51));
	U376 : AND3 port map(A1 => carry(48), A2 => p(48), A3 => p(49), Z => net_159);
	U377 : AND2 port map(A1 => g(48), A2 => p(49), Z => net_160);
	U378 : OR3 port map(A1 => net_159, A2 => net_160, A3 => g(49), Z => carry(50));
	U379 : AND2 port map(A1 => carry(48), A2 => p(48), Z => net_161);
	U380 : OR2 port map(A1 => net_161, A2 => g(48), Z => carry(49));
	U381 : AND4 port map(A1 => carry(52), A2 => p(52), A3 => p(53), A4 => p(54), Z => net_162);
	U382 : AND3 port map(A1 => g(52), A2 => p(53), A3 => p(54), Z => net_163);
	U383 : AND2 port map(A1 => g(53), A2 => p(54), Z => net_164);
	U384 : OR4 port map(A1 => net_162, A2 => net_163, A3 => net_164, A4 => g(54), Z => carry(55));
	U385 : AND3 port map(A1 => carry(52), A2 => p(52), A3 => p(53), Z => net_165);
	U386 : AND2 port map(A1 => g(52), A2 => p(53), Z => net_166);
	U387 : OR3 port map(A1 => net_165, A2 => net_166, A3 => g(53), Z => carry(54));
	U388 : AND2 port map(A1 => carry(52), A2 => p(52), Z => net_167);
	U389 : OR2 port map(A1 => net_167, A2 => g(52), Z => carry(53));
	U390 : AND4 port map(A1 => carry(56), A2 => p(56), A3 => p(57), A4 => p(58), Z => net_168);
	U391 : AND3 port map(A1 => g(56), A2 => p(57), A3 => p(58), Z => net_169);
	U392 : AND2 port map(A1 => g(57), A2 => p(58), Z => net_170);
	U393 : OR4 port map(A1 => net_168, A2 => net_169, A3 => net_170, A4 => g(58), Z => carry(59));
	U394 : AND3 port map(A1 => carry(56), A2 => p(56), A3 => p(57), Z => net_171);
	U395 : AND2 port map(A1 => g(56), A2 => p(57), Z => net_172);
	U396 : OR3 port map(A1 => net_171, A2 => net_172, A3 => g(57), Z => carry(58));
	U397 : AND2 port map(A1 => carry(56), A2 => p(56), Z => net_173);
	U398 : OR2 port map(A1 => net_173, A2 => g(56), Z => carry(57));
	U399 : AND4 port map(A1 => carry(60), A2 => p(60), A3 => p(61), A4 => p(62), Z => net_174);
	U400 : AND3 port map(A1 => g(60), A2 => p(61), A3 => p(62), Z => net_175);
	U401 : AND2 port map(A1 => g(61), A2 => p(62), Z => net_176);
	U402 : OR4 port map(A1 => net_174, A2 => net_175, A3 => net_176, A4 => g(62), Z => carry(63));
	U403 : AND3 port map(A1 => carry(60), A2 => p(60), A3 => p(61), Z => net_177);
	U404 : AND2 port map(A1 => g(60), A2 => p(61), Z => net_178);
	U405 : OR3 port map(A1 => net_177, A2 => net_178, A3 => g(61), Z => carry(62));
	U406 : AND2 port map(A1 => carry(60), A2 => p(60), Z => net_179);
	U407 : OR2 port map(A1 => net_179, A2 => g(60), Z => carry(61));
	U408 : XOR2 port map(A1 => carry(0), A2 => p(0), Z => sum(0));
	U409 : XOR2 port map(A1 => carry(1), A2 => p(1), Z => sum(1));
	U410 : XOR2 port map(A1 => carry(2), A2 => p(2), Z => sum(2));
	U411 : XOR2 port map(A1 => carry(3), A2 => p(3), Z => sum(3));
	U412 : XOR2 port map(A1 => carry(4), A2 => p(4), Z => sum(4));
	U413 : XOR2 port map(A1 => carry(5), A2 => p(5), Z => sum(5));
	U414 : XOR2 port map(A1 => carry(6), A2 => p(6), Z => sum(6));
	U415 : XOR2 port map(A1 => carry(7), A2 => p(7), Z => sum(7));
	U416 : XOR2 port map(A1 => carry(8), A2 => p(8), Z => sum(8));
	U417 : XOR2 port map(A1 => carry(9), A2 => p(9), Z => sum(9));
	U418 : XOR2 port map(A1 => carry(10), A2 => p(10), Z => sum(10));
	U419 : XOR2 port map(A1 => carry(11), A2 => p(11), Z => sum(11));
	U420 : XOR2 port map(A1 => carry(12), A2 => p(12), Z => sum(12));
	U421 : XOR2 port map(A1 => carry(13), A2 => p(13), Z => sum(13));
	U422 : XOR2 port map(A1 => carry(14), A2 => p(14), Z => sum(14));
	U423 : XOR2 port map(A1 => carry(15), A2 => p(15), Z => sum(15));
	U424 : XOR2 port map(A1 => carry(16), A2 => p(16), Z => sum(16));
	U425 : XOR2 port map(A1 => carry(17), A2 => p(17), Z => sum(17));
	U426 : XOR2 port map(A1 => carry(18), A2 => p(18), Z => sum(18));
	U427 : XOR2 port map(A1 => carry(19), A2 => p(19), Z => sum(19));
	U428 : XOR2 port map(A1 => carry(20), A2 => p(20), Z => sum(20));
	U429 : XOR2 port map(A1 => carry(21), A2 => p(21), Z => sum(21));
	U430 : XOR2 port map(A1 => carry(22), A2 => p(22), Z => sum(22));
	U431 : XOR2 port map(A1 => carry(23), A2 => p(23), Z => sum(23));
	U432 : XOR2 port map(A1 => carry(24), A2 => p(24), Z => sum(24));
	U433 : XOR2 port map(A1 => carry(25), A2 => p(25), Z => sum(25));
	U434 : XOR2 port map(A1 => carry(26), A2 => p(26), Z => sum(26));
	U435 : XOR2 port map(A1 => carry(27), A2 => p(27), Z => sum(27));
	U436 : XOR2 port map(A1 => carry(28), A2 => p(28), Z => sum(28));
	U437 : XOR2 port map(A1 => carry(29), A2 => p(29), Z => sum(29));
	U438 : XOR2 port map(A1 => carry(30), A2 => p(30), Z => sum(30));
	U439 : XOR2 port map(A1 => carry(31), A2 => p(31), Z => sum(31));
	U440 : XOR2 port map(A1 => carry(32), A2 => p(32), Z => sum(32));
	U441 : XOR2 port map(A1 => carry(33), A2 => p(33), Z => sum(33));
	U442 : XOR2 port map(A1 => carry(34), A2 => p(34), Z => sum(34));
	U443 : XOR2 port map(A1 => carry(35), A2 => p(35), Z => sum(35));
	U444 : XOR2 port map(A1 => carry(36), A2 => p(36), Z => sum(36));
	U445 : XOR2 port map(A1 => carry(37), A2 => p(37), Z => sum(37));
	U446 : XOR2 port map(A1 => carry(38), A2 => p(38), Z => sum(38));
	U447 : XOR2 port map(A1 => carry(39), A2 => p(39), Z => sum(39));
	U448 : XOR2 port map(A1 => carry(40), A2 => p(40), Z => sum(40));
	U449 : XOR2 port map(A1 => carry(41), A2 => p(41), Z => sum(41));
	U450 : XOR2 port map(A1 => carry(42), A2 => p(42), Z => sum(42));
	U451 : XOR2 port map(A1 => carry(43), A2 => p(43), Z => sum(43));
	U452 : XOR2 port map(A1 => carry(44), A2 => p(44), Z => sum(44));
	U453 : XOR2 port map(A1 => carry(45), A2 => p(45), Z => sum(45));
	U454 : XOR2 port map(A1 => carry(46), A2 => p(46), Z => sum(46));
	U455 : XOR2 port map(A1 => carry(47), A2 => p(47), Z => sum(47));
	U456 : XOR2 port map(A1 => carry(48), A2 => p(48), Z => sum(48));
	U457 : XOR2 port map(A1 => carry(49), A2 => p(49), Z => sum(49));
	U458 : XOR2 port map(A1 => carry(50), A2 => p(50), Z => sum(50));
	U459 : XOR2 port map(A1 => carry(51), A2 => p(51), Z => sum(51));
	U460 : XOR2 port map(A1 => carry(52), A2 => p(52), Z => sum(52));
	U461 : XOR2 port map(A1 => carry(53), A2 => p(53), Z => sum(53));
	U462 : XOR2 port map(A1 => carry(54), A2 => p(54), Z => sum(54));
	U463 : XOR2 port map(A1 => carry(55), A2 => p(55), Z => sum(55));
	U464 : XOR2 port map(A1 => carry(56), A2 => p(56), Z => sum(56));
	U465 : XOR2 port map(A1 => carry(57), A2 => p(57), Z => sum(57));
	U466 : XOR2 port map(A1 => carry(58), A2 => p(58), Z => sum(58));
	U467 : XOR2 port map(A1 => carry(59), A2 => p(59), Z => sum(59));
	U468 : XOR2 port map(A1 => carry(60), A2 => p(60), Z => sum(60));
	U469 : XOR2 port map(A1 => carry(61), A2 => p(61), Z => sum(61));
	U470 : XOR2 port map(A1 => carry(62), A2 => p(62), Z => sum(62));
	U471 : XOR2 port map(A1 => carry(63), A2 => p(63), Z => sum(63));
end struct;
